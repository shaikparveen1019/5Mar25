file2
Hello
